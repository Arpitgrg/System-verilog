`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 15.11.2023 15:55:12
// Design Name: 
// Module Name: mux_21
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux_21(
                    input a_in,
                    input b_in,
                    input sel,
                    output logic y_out);
always@*
begin

        case(sel)
        1'b0 :y_out= a_in;
        1'b1 :y_out=b_in;
        endcase
end                   
endmodule
